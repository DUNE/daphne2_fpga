-- st40_top.vhd
-- DAPHNE core logic, top level, self triggered mode sender
-- all 40 AFE channels -> one output link to DAQ
-- 
-- Jamieson Olsen <jamieson@fnal.gov>

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

use work.daphne2_package.all;

entity st40_top is
generic( link_id: std_logic_vector(5 downto 0)  := "000000" ); -- this is the OUTPUT link ID that goes into the header
port(
    reset: in std_logic;

    adhoc: in std_logic_vector(7 downto 0); -- user defined command for adhoc trigger
    threshold: in std_logic_vector(13 downto 0); -- user defined threshold relative to avg baseline
    ti_trigger: in std_logic_vector(7 downto 0); -------------------------
    ti_trigger_stbr: in std_logic;  -------------------------
    trig_rst_count: in std_logic;
    slot_id: in std_logic_vector(3 downto 0);
    crate_id: in std_logic_vector(9 downto 0);
    detector_id: in std_logic_vector(5 downto 0);
    version_id: in std_logic_vector(5 downto 0);
    enable: in std_logic_vector(39 downto 0);

    aclk: in std_logic; -- AFE clock 62.500 MHz
    timestamp: in std_logic_vector(63 downto 0);
	afe_dat: in array_5x9x14_type; -- ALL AFE channels feed into this module

    fclk: in std_logic; -- transmit clock to FELIX 120.237 MHz 
    dout: out std_logic_vector(31 downto 0);
    kout: out std_logic_vector(3 downto 0);
    Rcount_addr: in std_logic_vector(6 downto 0);
    Rcount: out std_logic_vector(63 downto 0)
    
);
end st40_top;

architecture st40_top_arch of st40_top is
 
    type state_type is (rst, scan, dump);
    signal state: state_type;

    signal sela: integer range 0 to 4;
    signal selc: integer range 0 to 7;
    signal sela_rden: integer range 0 to 4;
    signal selc_rden: integer range 0 to 7;
    signal fifo_ae: array_5x8_type;
    signal fifo_rden: array_5x8_type;
    signal fifo_ready: std_logic;
    signal fifo_do: array_5x8x32_type;
    signal fifo_ko: array_5x8x4_type;
    signal d, dout_reg: std_logic_vector(31 downto 0);
    signal k, kout_reg: std_logic_vector( 3 downto 0);
    signal packet_size_counter: integer range 0 to 467;
    signal trigcount: array_5x8x64_type;
    signal packcount: array_5x8x64_type;
    signal sendCount: unsigned(63 downto 0) := (others => '0');

    component stc is
    generic( link_id: std_logic_vector(5 downto 0) := "000000"; ch_id: std_logic_vector(5 downto 0) := "000000" );
    port(
        reset: in std_logic;

        adhoc: in std_logic_vector(7 downto 0);
        threshold: std_logic_vector(13 downto 0);
        slot_id: std_logic_vector(3 downto 0);
        crate_id: std_logic_vector(9 downto 0);
        detector_id: std_logic_vector(5 downto 0);
        version_id: std_logic_vector(5 downto 0);
        enable: std_logic;

        aclk: in std_logic; -- AFE clock 62.500 MHz
        timestamp: in std_logic_vector(63 downto 0);
    	ti_trigger: in std_logic_vector(7 downto 0); -------------------------
        ti_trigger_stbr: in std_logic;  -------------------------
        trig_rst_count: in std_logic;
        afe_dat: in std_logic_vector(13 downto 0);
        fclk: in std_logic; -- transmit clock to FELIX 120.237 MHz 
        fifo_rden: in std_logic;
        fifo_ae: out std_logic;
        fifo_do: out std_logic_vector(31 downto 0);
        fifo_ko: out std_logic_vector( 3 downto 0);
        Tcount: out std_logic_vector(63 downto 0);
        Pcount: out std_logic_vector(63 downto 0)
      );
    end component;

begin

    -- make 40 STC machines to monitor 40 AFE channels

    gen_stc_a: for a in 4 downto 0 generate
        gen_stc_c: for c in 7 downto 0 generate

            stc_inst: stc 
            generic map( link_id => link_id, ch_id => std_logic_vector(to_unsigned(10*a+c,6)) ) 
            port map(
                reset => reset,
    
                adhoc => adhoc,
                threshold => threshold,
                ti_trigger => ti_trigger, -------------------------
                ti_trigger_stbr => ti_trigger_stbr,  -------------------------
                trig_rst_count => trig_rst_count,
                slot_id => slot_id,
                crate_id => crate_id,
                detector_id => detector_id,
                version_id => version_id,
                enable => enable(8*a+c),
    
                aclk => aclk,
                timestamp => timestamp,
            	afe_dat => afe_dat(a)(c),
                fclk => fclk,
                fifo_rden => fifo_rden(a)(c),
                fifo_ae => fifo_ae(a)(c),
                fifo_do => fifo_do(a)(c),
                fifo_ko => fifo_ko(a)(c),
                Tcount => trigcount(a)(c),
                Pcount => packcount(a)(c)
              );

    end generate gen_stc_c;
    end generate gen_stc_a;

    -- fifo read enable and fifo flag selection

--    fifo_ready <= '1' when (sel_reg="000000" and fifo_ae(0)='1') else 
--                  '1' when (sel_reg="000001" and fifo_ae(1)='1') else 
--                  '1' when (sel_reg="000010" and fifo_ae(2)='1') else 
--                  '1' when (sel_reg="000011" and fifo_ae(3)='1') else 
--                  '1' when (sel_reg="000100" and fifo_ae(4)='1') else 
--                  '1' when (sel_reg="000101" and fifo_ae(5)='1') else 
--                  '1' when (sel_reg="000110" and fifo_ae(6)='1') else 
--                  '1' when (sel_reg="000111" and fifo_ae(7)='1') else 
--                  '1' when (sel_reg="001000" and fifo_ae(8)='1') else 
--                  '1' when (sel_reg="001001" and fifo_ae(9)='1') else 
--                  '0';

    -- sel_reg is a straight 6 bit register, but it is encoded with values 0-7, 10-17, 20-27, 30-37, 40-47
    -- there are gaps, so be careful when incrementing and looping...

    fifo_ready_proc: process(sela, selc, fifo_ae)
    begin
        fifo_ready <= '0'; -- default
        loop_a: for a in 4 downto 0 loop
            loop_c: for c in 7 downto 0 loop
                if (sela=a and selc=c and fifo_ae(a)(c)='1') then
                    fifo_ready <= '1';
                end if;
            end loop loop_c;
        end loop loop_a;
    end process fifo_ready_proc;

    gen_rden_a: for a in 4 downto 0 generate
        gen_rden_c: for c in 7 downto 0 generate
            fifo_rden(a)(c) <= '1' when (sela_rden=a and selc_rden=c and state=dump) else '0';
        end generate gen_rden_c;
    end generate gen_rden_a;

    -- FSM scans all STC machines in round robin manner, looking for a FIFO almost empty "fifo_ae" flag set. when it finds
    -- this, it reads one complete frame from that machine, then sends a few idles, then returns to scanning again.

    fsm_proc: process(fclk)
    begin
        if rising_edge(fclk) then
            if (reset='1' or trig_rst_count='1') then 
                state <= rst;
                sendCount <= (others => '0');
            else
                case(state) is

                    when rst =>
                        sela <= 0;
                        selc <= 0;
                        state <= scan;

                    when scan => 
                        if (trig_rst_count = '1') then
                            sendCount <= (others => '0');
                        end if;
                        if (fifo_ready='1') then
                            state <= dump;
                            sela_rden <= sela; 
                            selc_rden <= selc; 
                        else
                            state <= scan;
                        end if;
                        if (selc=7) then
                            if (sela=4) then -- loop around when sel = 4 7
                                sela <= 0;
                                selc <= 0;
                            else
                                sela <= sela + 1;
                                selc <= 0;
                            end if;
                        else
                            selc <= selc + 1;
                        end if;
                        packet_size_counter <= 0;
                    when dump =>
                        if (trig_rst_count = '1') then
                            sendCount <= (others => '0');
                        end if;
                        if ((k="0001" and d(7 downto 0)=X"DC") or packet_size_counter=467) then -- this the EOF word, done reading from this STC
                            state <= scan;
                            sendCount <= sendCount + 1;
                        else
                            state <= dump; -- in this state I can continue to search for the next fifo_ready_flag
                            packet_size_counter <= packet_size_counter + 1;
                            if (fifo_ready='0') then
                                if (selc=7) then
                                    if (sela=4) then -- loop around when sel = 4 7
                                        sela <= 0;
                                        selc <= 0;
                                    else
                                        sela <= sela + 1;
                                        selc <= 0;
                                    end if;
                                else
                                    selc <= selc + 1;
                                end if;   
                            end if;
                        end if;
                    when others => 
                        state <= rst;
                end case;
            end if;
        end if;
    end process fsm_proc;

    -- output muxes
     
--    d <= fifo_do(0) when (sel_reg="000000" and state=dump) else
--         fifo_do(1) when (sel_reg="000001" and state=dump) else
--         fifo_do(2) when (sel_reg="000010" and state=dump) else
--         fifo_do(3) when (sel_reg="000011" and state=dump) else
--         fifo_do(4) when (sel_reg="000100" and state=dump) else
--         fifo_do(5) when (sel_reg="000101" and state=dump) else
--         fifo_do(6) when (sel_reg="000110" and state=dump) else
--         fifo_do(7) when (sel_reg="000111" and state=dump) else
--         fifo_do(8) when (sel_reg="001000" and state=dump) else
--         fifo_do(9) when (sel_reg="001001" and state=dump) else
--         X"000000BC"; -- idle word
--
--    k <= fifo_ko(0) when (sel_reg="000000" and state=dump) else
--         fifo_ko(1) when (sel_reg="000001" and state=dump) else
--         fifo_ko(2) when (sel_reg="000010" and state=dump) else
--         fifo_ko(3) when (sel_reg="000011" and state=dump) else
--         fifo_ko(4) when (sel_reg="000100" and state=dump) else
--         fifo_ko(5) when (sel_reg="000101" and state=dump) else
--         fifo_ko(6) when (sel_reg="000110" and state=dump) else
--         fifo_ko(7) when (sel_reg="000111" and state=dump) else
--         fifo_ko(8) when (sel_reg="001000" and state=dump) else
--         fifo_ko(9) when (sel_reg="001001" and state=dump) else
--         "0001"; -- idle word

    outmux_proc: process(fifo_do, fifo_ko, sela_rden, selc_rden, state, packet_size_counter)
    begin
        d <= X"000000BC"; -- default
        k <= "0001"; -- default
        loop_a: for a in 4 downto 0 loop
        loop_c: for c in 7 downto 0 loop
            if ( sela_rden=a and selc_rden=c and state=dump ) then
                if (packet_size_counter=467 and fifo_ko(a)(c) /= "0001" and fifo_do(a)(c) /= X"DC") then
                    d <= X"011223DC";     
                    k <= "0001";
                else
                    d <= fifo_do(a)(c);
                    k <= fifo_ko(a)(c);
                end if;
            end if;
        end loop loop_c;
        end loop loop_a;
    end process outmux_proc;

    -- register the outputs

    outreg_proc: process(fclk)
    begin
        if rising_edge(fclk) then
            dout_reg <= d;
            kout_reg <= k;
        end if;
    end process outreg_proc;

    dout <= dout_reg;
    kout <= kout_reg;
    
    rcount_mux_proc: process(fclk)
    begin 
        if rising_edge(fclk) then
            case Rcount_addr is
                when std_logic_vector(to_unsigned(0,7)) =>
                    Rcount <= trigcount(0)(0);
                when std_logic_vector(to_unsigned(1,7)) =>
                    Rcount <= trigcount(0)(1);
                when std_logic_vector(to_unsigned(2,7)) =>
                    Rcount <= trigcount(0)(2);
                when std_logic_vector(to_unsigned(3,7)) =>
                    Rcount <= trigcount(0)(3);
                when std_logic_vector(to_unsigned(4,7)) =>
                    Rcount <= trigcount(0)(4);
                when std_logic_vector(to_unsigned(5,7)) =>
                    Rcount <= trigcount(0)(5);
                when std_logic_vector(to_unsigned(6,7)) =>
                    Rcount <= trigcount(0)(6);
                when std_logic_vector(to_unsigned(7,7)) =>
                    Rcount <= trigcount(0)(7);
                when std_logic_vector(to_unsigned(8,7)) =>
                    Rcount <= trigcount(1)(0);
                when std_logic_vector(to_unsigned(9,7)) =>
                    Rcount <= trigcount(1)(1);
                when std_logic_vector(to_unsigned(10,7)) =>
                    Rcount <= trigcount(1)(2);
                when std_logic_vector(to_unsigned(11,7)) =>
                    Rcount <= trigcount(1)(3);
                when std_logic_vector(to_unsigned(12,7)) =>
                    Rcount <= trigcount(1)(4);
                when std_logic_vector(to_unsigned(13,7)) =>
                    Rcount <= trigcount(1)(5);
                when std_logic_vector(to_unsigned(14,7)) =>
                    Rcount <= trigcount(1)(6);
                when std_logic_vector(to_unsigned(15,7)) =>
                    Rcount <= trigcount(1)(7);
                when std_logic_vector(to_unsigned(16,7)) =>
                    Rcount <= trigcount(2)(0);
                when std_logic_vector(to_unsigned(17,7)) =>
                    Rcount <= trigcount(2)(1);
                when std_logic_vector(to_unsigned(18,7)) =>
                    Rcount <= trigcount(2)(2);
                when std_logic_vector(to_unsigned(19,7)) =>
                    Rcount <= trigcount(2)(3);
                when std_logic_vector(to_unsigned(20,7)) =>
                    Rcount <= trigcount(2)(4);
                when std_logic_vector(to_unsigned(21,7)) =>
                    Rcount <= trigcount(2)(5);
                when std_logic_vector(to_unsigned(22,7)) =>
                    Rcount <= trigcount(2)(6);
                when std_logic_vector(to_unsigned(23,7)) =>
                    Rcount <= trigcount(2)(7);
                when std_logic_vector(to_unsigned(24,7)) =>
                    Rcount <= trigcount(3)(0);
                when std_logic_vector(to_unsigned(25,7)) =>
                    Rcount <= trigcount(3)(1);
                when std_logic_vector(to_unsigned(26,7)) =>
                    Rcount <= trigcount(3)(2);
                when std_logic_vector(to_unsigned(27,7)) =>
                    Rcount <= trigcount(3)(3);
                when std_logic_vector(to_unsigned(28,7)) =>
                    Rcount <= trigcount(3)(4);
                when std_logic_vector(to_unsigned(29,7)) =>
                    Rcount <= trigcount(3)(5);
                when std_logic_vector(to_unsigned(30,7)) =>
                    Rcount <= trigcount(3)(6);
                when std_logic_vector(to_unsigned(31,7)) =>
                    Rcount <= trigcount(3)(7);
                when std_logic_vector(to_unsigned(32,7)) =>
                    Rcount <= trigcount(4)(0);
                when std_logic_vector(to_unsigned(33,7)) =>
                    Rcount <= trigcount(4)(1);
                when std_logic_vector(to_unsigned(34,7)) =>
                    Rcount <= trigcount(4)(2);
                when std_logic_vector(to_unsigned(35,7)) =>
                    Rcount <= trigcount(4)(3);
                when std_logic_vector(to_unsigned(36,7)) =>
                    Rcount <= trigcount(4)(4);
                when std_logic_vector(to_unsigned(37,7)) =>
                    Rcount <= trigcount(4)(5);
                when std_logic_vector(to_unsigned(38,7)) =>
                    Rcount <= trigcount(4)(6);
                when std_logic_vector(to_unsigned(39,7)) =>
                    Rcount <= trigcount(4)(7);
                when std_logic_vector(to_unsigned(40,7)) =>
                    Rcount <= packcount(0)(0);
                when std_logic_vector(to_unsigned(41,7)) =>
                    Rcount <= packcount(0)(1);
                when std_logic_vector(to_unsigned(42,7)) =>
                    Rcount <= packcount(0)(2);
                when std_logic_vector(to_unsigned(43,7)) =>
                    Rcount <= packcount(0)(3);
                when std_logic_vector(to_unsigned(44,7)) =>
                    Rcount <= packcount(0)(4);
                when std_logic_vector(to_unsigned(45,7)) =>
                    Rcount <= packcount(0)(5);
                when std_logic_vector(to_unsigned(46,7)) =>
                    Rcount <= packcount(0)(6);
                when std_logic_vector(to_unsigned(47,7)) =>
                    Rcount <= packcount(0)(7);
                when std_logic_vector(to_unsigned(48,7)) =>
                    Rcount <= packcount(1)(0);
                when std_logic_vector(to_unsigned(49,7)) =>
                    Rcount <= packcount(1)(1);
                when std_logic_vector(to_unsigned(50,7)) =>
                    Rcount <= packcount(1)(2);
                when std_logic_vector(to_unsigned(51,7)) =>
                    Rcount <= packcount(1)(3);
                when std_logic_vector(to_unsigned(52,7)) =>
                    Rcount <= packcount(1)(4);
                when std_logic_vector(to_unsigned(53,7)) =>
                    Rcount <= packcount(1)(5);
                when std_logic_vector(to_unsigned(54,7)) =>
                    Rcount <= packcount(1)(6);
                when std_logic_vector(to_unsigned(55,7)) =>
                    Rcount <= packcount(1)(7);
                when std_logic_vector(to_unsigned(56,7)) =>
                    Rcount <= packcount(2)(0);
                when std_logic_vector(to_unsigned(57,7)) =>
                    Rcount <= packcount(2)(1);
                when std_logic_vector(to_unsigned(58,7)) =>
                    Rcount <= packcount(2)(2);
                when std_logic_vector(to_unsigned(59,7)) =>
                    Rcount <= packcount(2)(3);
                when std_logic_vector(to_unsigned(60,7)) =>
                    Rcount <= packcount(2)(4);
                when std_logic_vector(to_unsigned(61,7)) =>
                    Rcount <= packcount(2)(5);
                when std_logic_vector(to_unsigned(62,7)) =>
                    Rcount <= packcount(2)(6);
                when std_logic_vector(to_unsigned(63,7)) =>
                    Rcount <= packcount(2)(7);
                when std_logic_vector(to_unsigned(64,7)) =>
                    Rcount <= packcount(3)(0);
                when std_logic_vector(to_unsigned(65,7)) =>
                    Rcount <= packcount(3)(1);
                when std_logic_vector(to_unsigned(66,7)) =>
                    Rcount <= packcount(3)(2);
                when std_logic_vector(to_unsigned(67,7)) =>
                    Rcount <= packcount(3)(3);
                when std_logic_vector(to_unsigned(68,7)) =>
                    Rcount <= packcount(3)(4);
                when std_logic_vector(to_unsigned(69,7)) =>
                    Rcount <= packcount(3)(5);
                when std_logic_vector(to_unsigned(70,7)) =>
                    Rcount <= packcount(3)(6);
                when std_logic_vector(to_unsigned(71,7)) =>
                    Rcount <= packcount(3)(7);
                when std_logic_vector(to_unsigned(72,7)) =>
                    Rcount <= packcount(4)(0);
                when std_logic_vector(to_unsigned(73,7)) =>
                    Rcount <= packcount(4)(1);
                when std_logic_vector(to_unsigned(74,7)) =>
                    Rcount <= packcount(4)(2);
                when std_logic_vector(to_unsigned(75,7)) =>
                    Rcount <= packcount(4)(3);
                when std_logic_vector(to_unsigned(76,7)) =>
                    Rcount <= packcount(4)(4);
                when std_logic_vector(to_unsigned(77,7)) =>
                    Rcount <= packcount(4)(5);
                when std_logic_vector(to_unsigned(78,7)) =>
                    Rcount <= packcount(4)(6);
                when std_logic_vector(to_unsigned(79,7)) =>
                    Rcount <= packcount(4)(7);
                when std_logic_vector(to_unsigned(80,7)) =>
                    Rcount <= std_logic_vector(sendCount);
                when others => 
                    Rcount <= (others => '1');
            end case;
        end if;
    end process rcount_mux_proc;

end st40_top_arch;